//Verilog HDL for "Lib6710_02", "TIEHI" "behavioral"


module TIEHI ( Y );

  output Y;

  assign Y = 1'b1;

endmodule

