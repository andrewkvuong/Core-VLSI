//Verilog HDL for "Lib6710_02", "TIELO" "behavioral"


module TIELO ( Y );

  output Y;

  assign Y = 1'b0;

endmodule
